library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity ROM is
 port(
 address : in std_logic_vector(3 downto 0);
 dout : out std_logic_vector(3 downto 0)
 );
end entity ROM;
architecture RTL of ROM is
 type MEMORY_16_4 is array (0 to 15) of std_logic_vector(3 downto 0);
 constant ROM_16_4 : MEMORY_16_4 := (
 x"0",
 x"1",
 x"2",
 x"3",
 x"4",
 x"5",
 x"6",
 x"7",
 x"8",
 x"9",
 x"a",
 x"b",
 x"c",
 x"d",
 x"e",
 x"f"
 );
begin
 main : process(address)
 begin
 dout <= ROM_16_4(to_integer(unsigned(address)));
 end process main;
end architecture RTL;